module practica2
(
	input clk,
	input reset, 
	input Enable,
	
	output tiempo
);




endmodule 