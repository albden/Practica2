module practica2
(
	input clk,
	input reset, 
	input Enable,
	input start,
	
	output tiempo
);




endmodule 
