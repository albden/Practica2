module practica2
(
	input clk,
	input reset, 
	input Enable,
	input start,
	input entrada_A,
	input entrada_B,
		
	output tiempo,
	output product,
	output Clk
);




endmodule 
